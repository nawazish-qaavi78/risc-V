
// datapath.v
module datapath (
    input         clk, reset,
    input [1:0]   ResultSrc, PCSrc,
    input         ALUSrc,
    input         RegWrite, 
    input [2:0]   ImmSrc,
    input [3:0]   ALUControl,
    output [3:0]       flags,
    output [31:0] PC,
    input  [31:0] Instr,
    output [31:0] Mem_WrAddr, Mem_WrData,
    input  [31:0] ReadData,
    output [31:0] Result
);

wire [31:0] PCNext, PCPlus4, PCTarget, UOut;
wire [31:0] ImmExt, SrcA, SrcB, WriteData, ALUResult;
wire [31:0] PCadd_result;


// next PC logic
reset_ff #(32) pcreg(clk, reset, PCNext, PC);

adder 			pcadd(PC, (PCSrc[0]?32'd4:ImmExt), PCadd_result);
assign PCPlus4 = (PCSrc[0] == 0) ? PCadd_result : 32'b0;
assign PCTarget = (PCSrc[0] == 1) ? PCadd_result : 32'b0;


mux3 #(32)     pcmux(PCPlus4, PCTarget, ALUResult, PCSrc, PCNext);

mux2 #(32)		umux(PCTarget, ImmExt, Instr[5], UOut);

// register file logic
reg_file       rf (clk, RegWrite, Instr[19:15], Instr[24:20], Instr[11:7], Result, SrcA, WriteData);
imm_extend     ext (Instr[31:7], ImmSrc, ImmExt);

// ALU logic
mux2 #(32)     srcbmux(WriteData, ImmExt, ALUSrc, SrcB);
alu            alu (SrcA, SrcB, ALUControl, ALUResult, flags);
mux4 #(32)     resultmux(ALUResult, ReadData, PCPlus4, UOut, ResultSrc, Result);


assign Mem_WrData = WriteData;
assign Mem_WrAddr = ALUResult;

endmodule

